// Verilog
// woStLN
// Ninputs 2
// Noutputs 1
// NtotalGates 25
// BUF1 1
// NAND2 20
// NAND3 4

module  woStLN (N11,N14,N90);

input N11,N14;

output N90;

wire N118,N119,N122,N123,N124,N125,N126,N218,N219,N222,
     N223,N224,N225,N226,N248,N249,N242,N243,N244,N245,
     N246,N250,N251,N252,N253,N254,N255,N256;

nand NAND2_1 (N126, N125, N124);
nand NAND2_2 (N125, N11, N123);
nand NAND2_3 (N124, N126, N14);
nand NAND3_4 (N123, N124, N125, N14);
nand NAND2_5 (N119, N118, N123);
nand NAND2_6 (N118, N119, N124);
nand NAND2_7 (N226, N225, N224);
nand NAND2_8 (N225, N118, N223);
nand NAND2_9 (N224, N226, N14);
nand NAND3_10 (N223, N224, N225, N14);
nand NAND2_11 (N219, N218, N223);
nand NAND2_12 (N218, N219, N224);
nand NAND2_13 (N246, N245, N244);
nand NAND2_14 (N245, N218, N243);
nand NAND2_15 (N244, N246, N14);
nand NAND3_16 (N243, N244, N245, N14);
nand NAND2_17 (N249, N248, N243);
nand NAND2_18 (N248, N249, N244);
nand NAND2_19 (N256, N255, N254);
nand NAND2_20 (N255, N248, N253);
nand NAND2_21 (N254, N256, N14);
nand NAND3_22 (N253, N254, N255, N14);
nand NAND2_23 (N251, N250, N253);
nand NAND2_24 (N250, N251, N254);
buf BUF_25 (N90, N250);

endmodule
